GC AULT                                 D�� D��               L1152                   @4��    @P�&�   D��D��              L1172                   @5�`   @P�    D��D��              L1498                   @���   @9	u@   D��D��              Taurus                  @�f`   @;���   D�� D��               b1498                   @���   @9	u@   D��D��              c778                    @3h?�   @7�`   D��D��              ON1                     @44�`   @?�     D��D��              L1641 T                 @$�O��r�       D�� D��               Pleiades                @Ǯ    @7s3@   D�� D��               s255  8                 @���   @2l    D�� D��               S255  8                 @���   @2l    D�� D��               OrionB                  @��    �����   D�� D��               RNO43                   @��   @)��    D�� D��               IRC+ LT                 @#�"    @+f`   D�� D��               RMon  8                 @mˠ   @!���   D�� D��               Ori18 T                 @/�������"""""D�� D��               DR21  T                 @4��`   @E�    D�� D��               MBM12 T                 @c�     �A333333D�� D��               G70+1.2                 @4
�@   @@�    D�� D��               S106 LT                 @4m�   @B�`�   D�� D��               W42   8                 @8ff`   �ə��   D�� D��               L111  T                 @[�             D�� D��               l134n T                 @/�wwwww�������D�� D��               ngc2264                 @��    @#�   D�� D��               outflow                 @5���   @G�Ӡ   D�� D��               CygX LT                 @T              D�� D��               KHW ULT                 @�q���       D�� D��               HH1-2 T                 @/��   ��"    D�� D��               IRASclouds              @�y�   �!�    D�� D��               BUBNEB                  @7N�@   @NuU�   D�� D��               L1228 T                 @4�w�   @SX��   D�� D��               ngc2071 AS              @�jAg        D�� D��               dr21  T                 @4��`   @E�    D�� D��               ngc1333                 @vT2��@?�%��YD�� D��               B5 1333                 @�]@   @@^�    D�� D��               MBM41 T                 @0�    @NuU`   D�� D��               OrionW                  @UU`   �33@   D�� D��               446-552                 @�`   �ww�   D�� D��               440-534                 @���-���UUUUUUD�� D��               NGC4449                 @(ۻ�   @F.��   D�� D��               hh83 84                 @�є#�������D�� D��               OriA LT                 @/��   ��"    D�� D��               S157 LT                 @7;��   @M���   D��D��              mbir LT                 @:�vT2@3ꪪ���D�� D��               BNKL LT                 @/�������"""""D�� D��               orib  T                 @��    �����   D�� D��               L134N T                 @/�w�   ����   D�� D��               MBM32 T                 @"��    @P�U`   D�� D��               NGP ULT                         @V�     D�� D��               l=110 T                 @[�             D�� D��               n7027 T                 @5�@   @E_�   D�� D��               MBM30 T                 @"΁�   @Q���   D�� D��               MBM27 T                 @!u   @R33@   D�� D��               irs5  1 AS              @�E��8@22J.�_D�� D�� �F�          SGRA LT                 @1�/�b���<������D�� D��               SGRA-LB                 @v�hr�!��?|�hsD�� D��               B5I4  5 AS              @�X�%��@@t_���,D�� D��               MBM41-LB                @V��>BZ�@C�*�1D�� D��               HPX ENS                 @��vT2@3>o����D�� D��               S159 LT                 @79�����@NuUUUUUD�� D��               M31 ULT                 ?�UU`   @De@   D�� D��               MBM26 T                 @ ��   @N[��   D�� D��               beichman                @�   @<f�   D�� D��               M31-2000                ?���,_��@D�"""""D�  D�                M31-XY                  ?�UUUUUU@DeC ��D�� D�� �J(�\     B5IRS4                  @�X�%��@@t_���,D�� D��               M3 A LT                 @+Tz�   @<�"    D�� D��               BG 32 T                 @#    @PZ��   D�� D��               MBM40 T                 @0#�    @5�3@   D�� D��               BGL1551                 @��[�@2      D�� D��               BG03  T                 @�33333@*      D�� D��               BG02  T                 @��[�@2      D�� D��               BGB301                  @�"""""@*ffffffD�� D��               BGB302                  @�33333@)�fffffD�� D��               BGB303                  @�33333@*�fffffD�� D��               BGB304                  @�33333@*ffffffD�� D��               BGB305                  @�33333@*ffffffD�� D��               BGB35                   @�UUUUU@"UUUUUUD�� D��               BGL15991                @�����@j�����D�� D��               BGL15992                @3����	@z�G�{D�� D��               BGs2471                 @t�I��J@5������D�� D��               BGs2472                 @t�I��J@5������D�� D��               BGs2551                 @��|�@2      D�� D��               BGs2552                 @��|�@2      D�� D��               BGs2553                 @��|�@2      D�� D��               BGs2554                 @���
=q@2      D�� D��               BGs2555                 @�T2��@2      D�� D��               BGmonfil                @UUUUUU@�i�6�D�� D��               BGMon1                  @������@*      D�� D��               BGMon2                  @������@%      D�� D��               BGMon3                  @������@%      D�� D��               BGMon4                  @������@$�     D�� D��               BGMon5                  @������@%�     D�� D��               BGL6661                 @2�UUUUU@/      D�� D��               BGL6662                 @2�UUUUU@.������D�� D��               BGL6663                 @2�UUUUU@/UUUUUUD�� D��               BGL6664                 @2�UUUUU@.UUUUUUD�� D��               BGL637                  @2�fffff@ @     D�� D��               BGfrog                  @2޸Q�@������D�� D��               BGL717                  @3&/�b��@1�UUUUUD�� D��               BGL7231                 @3Al�l@3�����D�� D��               BGL7232                 @3C���n@3�����D�� D��               BGL7233                 @3Al�l@3DDDDDDD�� D��               BGL7234                 @3Al�l@3n�����D�� D��               BGL6665                 @2�UUUUU@/������D�� D��               RaDec p3 S                              D�� D��                RADEC82  S                              D�� D��                IRS4 LT                 @�X�%��@@t_���,D�� D��               ISR4 LT                 @�X�%��@@t_���,D�� D��               CLOUD2                  @��m:�@9�UUUUUD�� D��               n1333 T                 @u0�   @?+��   D�� D��               c13135                  @1C�   @J���   D�� D��               c4055                   @a��   ����   D�� D��               c5270                   @�M@   @(r�   D�� D��               rosette                 @i�z�   ���    D�� D��               DR21(OH)                @4���   @E��   D�� D��               W49 ULT                 @3!��N�@"��5y�D�� D��               Orion A g               @/7�   ���    D�� D��               Orion_A g               @/7�   ���    D�� D��               