numpt
nver
nprc
nplc
onstk
nwts
locwt
ibsln
kuse
nstk
nlist
indx
isdum
numst
fwid
expch
refch
vlsr
exwid
wght
factt
time
pwrav
pwrer
rms
tmax
arerr
area
vcent
fwhm
fwerr
fpeak
fperr
ftmax
fterr
rmval
ra
dec
l
b
dra
ddec
dl
db
dx
dy
odra
oddec
epoch
vpeak
rsdm
freq
stak
nstkx
