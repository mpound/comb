	{"APPCAL",LOGICAL,APPCAL,48,10},
	{"BASELN",INT,BASELN,49,11},
	{"BITPIX",INT,BITPIX,1,0},
	{"BLANK",INT,BLANK,29,10},
	{"BSCALE",DOUBLE,BSCALE,30,10},
	{"BUNIT",STR,BUNIT,32,0},
	{"BZERO",DOUBLE,BZERO,31,10},
	{"CDELT1",DOUBLE,CDELT1,9,0},
	{"CDELT2",DOUBLE,CDELT2,14,0},
	{"CDELT3",DOUBLE,CDELT3,19,0},
	{"CDELT4",DOUBLE,CDELT4,24,0},
	{"CROTA1",DOUBLE,CROTA1,11,0},
	{"CROTA2",DOUBLE,CROTA2,16,0},
	{"CROTA3",DOUBLE,CROTA3,21,0},
	{"CROTA4",DOUBLE,CROTA4,26,0},
	{"CRPIX1",DOUBLE,CRPIX1,10,0},
	{"CRPIX2",DOUBLE,CRPIX2,15,0},
	{"CRPIX3",DOUBLE,CRPIX3,20,0},
	{"CRPIX4",DOUBLE,CRPIX4,25,0},
	{"CRVAL1",DOUBLE,CRVAL1,8,0},
	{"CRVAL2",DOUBLE,CRVAL2,13,0},
	{"CRVAL3",DOUBLE,CRVAL3,18,0},
	{"CRVAL4",DOUBLE,CRVAL4,23,0},
	{"CTYPE1",STR,CTYPE1,7,5},
	{"CTYPE2",STR,CTYPE2,12,6},
	{"CTYPE3",STR,CTYPE3,17,7},
	{"CTYPE4",STR,CTYPE4,22,8},
	{"DATAMAX",DOUBLE,DATAMAX,34,10},
	{"DATAMIN",DOUBLE,DATAMIN,33,10},
	{"DATE",STR,DATE,36,10},
	{"DATE-OBS",STR,DATEOBS,35,10},
	{"DELTAV",DOUBLE,DELTAV,46,11},
	{"END",LOGICAL,END,54,9},
	{"EPOCH",DOUBLE,EQUINOX,27,10},
	{"EQUINOX",DOUBLE,EQUINOX,28,10},
	{"IMAGEOP",IHISTORY,IMAGEOP,52,10},
	{"NAXIS",INT,NAXIS,2,0},
	{"NAXIS1",INT,NAXIS1,3,1},
	{"NAXIS2",INT,NAXIS2,4,2},
	{"NAXIS3",INT,NAXIS3,5,3},
	{"NAXIS4",INT,NAXIS4,6,4},
	{"OBJECT",STR,OBJECT,37,10},
	{"OBSTIME",DOUBLE,OBSTIME,44,11},
	{"PARAM",IHISTORY,PARAM,51,10},
	{"PROJTYPE",STR,PROJTYPE,47,10},
	{"RESTFREQ",DOUBLE,RESTFREQ,39,10},
	{"SCAN-NUM",DOUBLE,SCAN_NUM,40,11},
	{"SIMPLE",LOGICAL,SIMPLE,0,0},
	{"TELESCOP",STR,TELESCOP,38,10},
	{"TITLE",IHISTORY,TITLE,50,10},
	{"TSYS",DOUBLE,TSYS,45,11},
	{"USERHIST",IHISTORY,USERHIST,53,10},
	{"VELO",DOUBLE,VELO_LSR,43,11},
	{"VELO-LSR",DOUBLE,VELO_LSR,42,11},
	{"VLSR",DOUBLE,VELO_LSR,41,11}
